module bancoRegistradores(rst, clk, wrEn, addR1, addR2, addWr, dadoR1, dadoR2, dadoWr);
input clk, rst, wrEn;
input [2:0] addR1, addR2, addWr;
input [7:0] dadoWr;
output reg [7:0] dadoR1; 
output reg [7:0] dadoR2;

endmodule