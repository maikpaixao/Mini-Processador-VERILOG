module ula (portA, portB, op, resultado);
	input [7:0]portA; 
	input [7:0]portB; 
	input [2:0]op; 
	output reg [7:0]resultado; 
	
endmodule
